.title KiCad schematic
J1 __J1
J2 __J2
R6 /ENABLE Net-_J1-Pin_1_ 0
R7 GND Net-_U1-RT/CLK_ 43k
R4 SYS_DCIN /ENABLE 332k
R5 GND /ENABLE 56.2k
C9 GND Net-_U1-COMP_ 14p
R8 Net-_C8-Pad2_ Net-_U1-COMP_ 9k
U1 __U1
C7 GND Net-_U1-SS/TR_ 0.025u
C8 GND Net-_C8-Pad2_ 51.1n
C1 SYS_DCIN GND 22uF 2201010609TR
C5 +5V GND 100u
D1 __D1
L1 /SW +5V 10u
R2 +5V /FB 52k
R3 /FB GND 11k
C3 /SW /BOOT 0.1u
.end
